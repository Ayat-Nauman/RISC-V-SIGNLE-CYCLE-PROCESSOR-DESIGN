module decoder(
	input logic 
	);
